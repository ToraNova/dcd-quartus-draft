entity dcd_draft is
end entity;

architecture sim of dcd_draft is
begin

	process is
	begin
	--this is the main process
		report "Hello DCD!";
		wait;
	

	end process;
end architecture;
